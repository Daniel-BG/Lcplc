package constants is
	attribute KEEP: string;
	constant KEEP_DEFAULT: string := "TRUE";

	attribute USE_DSP48 : string;
	constant USE_DSP48_ARITH_OP: string := "YES";
end constants;

package body constants is

end constants;