----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.02.2019 09:19:13
-- Design Name: 
-- Module Name: binary_dequantizer - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.constants.all;

entity BINARY_DEQUANTIZER is
	Generic (
		--0 leaves it the same
		SHIFT		: integer := 0;
		DATA_WIDTH	: integer := 16;
		USER_WIDTH	: integer := 1
	);
	Port (
		clk, rst: std_logic;
		input_ready	: out std_logic;
		input_valid	: in  std_logic;
		input_data	: in  std_logic_vector(DATA_WIDTH - 1 downto 0);
		input_last  : in  std_logic := '0';
		input_user	: in  std_logic_vector(USER_WIDTH - 1 downto 0) := (others => '0');
		output_ready: in  std_logic;
		output_valid: out std_logic;
		output_data	: out std_logic_vector(DATA_WIDTH - 1 downto 0);
		output_last : out std_logic;
		output_user : out std_logic_vector(USER_WIDTH - 1 downto 0)
	);
end BINARY_DEQUANTIZER;

architecture Behavioral of BINARY_DEQUANTIZER is

	signal input_sign_extended: std_logic_vector(DATA_WIDTH downto 0);
	signal abs_val: std_logic_vector(DATA_WIDTH downto 0);
	
	signal shifted_up: std_logic_vector(DATA_WIDTH downto 0);

	signal pre_out: std_logic_vector(DATA_WIDTH downto 0);
	attribute KEEP of pre_out: signal is KEEP_DEFAULT;
	
begin

	
	--no segmentation done yet
	output_valid <= input_valid;
	input_ready  <= output_ready;
	output_last  <= input_last;
	output_user  <= input_user;

	input_sign_extended <= input_data(DATA_WIDTH - 1) & input_data;
	abs_val <= input_sign_extended when input_data(DATA_WIDTH - 1) = '0' else std_logic_vector(-signed(input_sign_extended));
	
	gen_zero_shift: if SHIFT = 0 generate
		shifted_up <= abs_val;
	end generate;
	gen_shift: if SHIFT > 0 generate
		shifted_up <= abs_val(DATA_WIDTH - SHIFT downto 0) & (SHIFT - 1 downto 0 => '0');
	end generate;
	
	pre_out <= shifted_up when input_data(DATA_WIDTH - 1) = '0' else std_logic_vector(-signed(shifted_up));
	output_data <= pre_out(DATA_WIDTH - 1 downto 0);

end Behavioral;
