`define GOLDEN_ROOT_DIR "C:/Users/Daniel/Repositorios/Lcplc/test_data/"
`define GOLDEN_EXT ".smpl"

`define GOLDEN_ALPHA		{`GOLDEN_ROOT_DIR, "alpha", 		`GOLDEN_EXT}
`define GOLDEN_ALPHAN		{`GOLDEN_ROOT_DIR, "alphan", 		`GOLDEN_EXT}
`define GOLDEN_ALPHAD		{`GOLDEN_ROOT_DIR, "alphad", 		`GOLDEN_EXT}
`define GOLDEN_X 			{`GOLDEN_ROOT_DIR, "x", 			`GOLDEN_EXT}
`define GOLDEN_XHAT 		{`GOLDEN_ROOT_DIR, "xhat", 			`GOLDEN_EXT}
`define GOLDEN_XMEAN 		{`GOLDEN_ROOT_DIR, "xmean", 		`GOLDEN_EXT}
`define GOLDEN_XHATMEAN 	{`GOLDEN_ROOT_DIR, "xhatmean", 		`GOLDEN_EXT}
`define GOLDEN_PREDICTION 	{`GOLDEN_ROOT_DIR, "prediction",	`GOLDEN_EXT}
