`define GOLDEN_ROOT_DIR "C:/Users/Daniel/Repositorios/Lcplc/test_data/"
`define GOLDEN_EXT ".smpl"

`define GOLDEN_X_FIRSTB			{`GOLDEN_ROOT_DIR, "x_firstband",			`GOLDEN_EXT}
`define GOLDEN_X_FIRSTB_LAST_R	{`GOLDEN_ROOT_DIR, "x_firstband_last_r",	`GOLDEN_EXT}
`define GOLDEN_X_FIRSTB_LAST_S	{`GOLDEN_ROOT_DIR, "x_firstband_last_s",	`GOLDEN_EXT}
`define GOLDEN_XTILDE_FIRSTB	{`GOLDEN_ROOT_DIR, "xtilde_firstband",		`GOLDEN_EXT}

`define GOLDEN_X_OTHERBANDS		{`GOLDEN_ROOT_DIR, "x_otherbands",			`GOLDEN_EXT}
`define GOLDEN_XHAT 			{`GOLDEN_ROOT_DIR, "xhat", 					`GOLDEN_EXT}
`define GOLDEN_XHAT_LAST_S 		{`GOLDEN_ROOT_DIR, "xhat_last_s", 			`GOLDEN_EXT}
`define GOLDEN_XMEAN 			{`GOLDEN_ROOT_DIR, "xmean", 				`GOLDEN_EXT}
`define GOLDEN_XHATMEAN 		{`GOLDEN_ROOT_DIR, "xhatmean", 				`GOLDEN_EXT}
`define GOLDEN_ALPHA			{`GOLDEN_ROOT_DIR, "alpha", 				`GOLDEN_EXT}

`define GOLDEN_XTILDE_OTHERBANDS{`GOLDEN_ROOT_DIR, "xtilde_otherbands",		`GOLDEN_EXT}
`define GOLDEN_XTILDE_O_LAST_S	{`GOLDEN_ROOT_DIR, "xtilde_others_last_s",	`GOLDEN_EXT}

`define GOLDEN_X 				{`GOLDEN_ROOT_DIR, "x", 					`GOLDEN_EXT}
`define GOLDEN_X_LAST_S			{`GOLDEN_ROOT_DIR, "x_Last_s",				`GOLDEN_EXT}
`define GOLDEN_X_LAST_B			{`GOLDEN_ROOT_DIR, "x_last_b",				`GOLDEN_EXT}
`define GOLDEN_X_LAST_I			{`GOLDEN_ROOT_DIR, "x_last_i",				`GOLDEN_EXT}

`define GOLDEN_XTILDE		 	{`GOLDEN_ROOT_DIR, "xtilde",				`GOLDEN_EXT}
`define GOLDEN_XTILDE_LAST_S 	{`GOLDEN_ROOT_DIR, "xtilde_last_s",			`GOLDEN_EXT}

`define GOLDEN_XHATRAW	 		{`GOLDEN_ROOT_DIR, "xhatraw",				`GOLDEN_EXT}
`define GOLDEN_XHATRAW_LAST_S	{`GOLDEN_ROOT_DIR, "xhatraw_last_s",		`GOLDEN_EXT}
`define GOLDEN_XHATRAW_LAST_B	{`GOLDEN_ROOT_DIR, "xhatraw_last_b",		`GOLDEN_EXT}

`define GOLDEN_DFLAG	 		{`GOLDEN_ROOT_DIR, "dflag",					`GOLDEN_EXT}

`define GOLDEN_MERR		 		{`GOLDEN_ROOT_DIR, "merr",					`GOLDEN_EXT}
`define GOLDEN_KJ		 		{`GOLDEN_ROOT_DIR, "kj",					`GOLDEN_EXT}





`define GOLDEN_ALPHAN		{`GOLDEN_ROOT_DIR, "alphan", 		`GOLDEN_EXT}
`define GOLDEN_ALPHAD		{`GOLDEN_ROOT_DIR, "alphad", 		`GOLDEN_EXT}

`define GOLDEN_PREDICTION 	{`GOLDEN_ROOT_DIR, "prediction",	`GOLDEN_EXT}

`define GOLDEN_EZG_INPUT    {`GOLDEN_ROOT_DIR, "egz_input",		`GOLDEN_EXT}
`define GOLDEN_EZG_CODE     {`GOLDEN_ROOT_DIR, "egz_code",		`GOLDEN_EXT}
`define GOLDEN_EZG_LENGTH   {`GOLDEN_ROOT_DIR, "egz_quant",		`GOLDEN_EXT}
`define GOLDEN_GC_INPUT		{`GOLDEN_ROOT_DIR, "gc_input", 		`GOLDEN_EXT}
`define GOLDEN_GC_PARAM		{`GOLDEN_ROOT_DIR, "gc_param", 		`GOLDEN_EXT}
`define GOLDEN_GC_CODE		{`GOLDEN_ROOT_DIR, "gc_code", 		`GOLDEN_EXT}
`define GOLDEN_GC_LENGTH	{`GOLDEN_ROOT_DIR, "gc_quant",		`GOLDEN_EXT}
`define GOLDEN_OUTPUT		{`GOLDEN_ROOT_DIR, "output",		`GOLDEN_EXT}