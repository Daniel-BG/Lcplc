package data_types is
    type array_of_integers is array(integer range <>) of integer;
end package;

package body data_types is

end data_types;