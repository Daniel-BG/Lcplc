package constants is
	attribute KEEP: string;
	constant KEEP_DEFAULT: string := "FALSE";
end constants;

package body constants is

end constants;